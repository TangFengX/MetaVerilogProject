module top(
    input a,b,clk,
    output c
);
    assign c=a&b;
    
endmodule


